module determinant2x2 (
    input [31:0] A_flat,  
    input clock,
    output reg [7:0] det,
    output reg done,
    output reg overflow_flag
);

  
endmodule