module alu_multiplication_module(
  input [199:0] A_flat,
  input [199:0] B_flat,
  output reg [199:0] C_flat,
  output reg overflow_flag,
  output reg done
);

endmodule

