module alu_scalar_module(
  input [199:0] A_flat,
  input [7:0] scalar,
  output reg [199:0] C_flat,
  output reg overflow_flag,
  output reg done
);


endmodule
